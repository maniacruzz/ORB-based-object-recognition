library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

package Amogh_pkg is

	
	-- Array types

	type vector_8bit is array(natural range <>) of std_logic_vector(8-1 downto 0);
	type int_vector_8bit is array(natural range <>) of integer range 0 to 255;
	type vector_23bit is array(natural range <>) of std_logic_vector(23-1 downto 0);


	--constant test : int_vector_8bit(1023 downto 0) := (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0);
	--constant test : int_vector_8bit(1023 downto 0) := (7,   3,  16,  15,  10,   9,  17,  24,  10,   7,   9,   6,  24,   8,  10,  17,  11,  18,  27,   8,  14,  13,   5,  20,  14,  22,  15,   5,  29,  10,  20,   1,  23,  20,  14,  19,  11,  15,  24,  18,  18,  19,  27,  27,   4,  32,  20,  15,  11,  20,  15,   9,  31,   1,  26,  13,  14,  22,  18,  19,  21,  21,  20,  28,  11,  19,  16,  20,  11,  25,   7,  19,  12,   5,   6,  22,  29,  21,  17,  17,  17,  19,  13,  20,  15,  27,  16,  25,  30,  20,   6,   7,  27,  22,  22,  16,  11,  15,   7,   7,  10,   7,  15,   7,  29,   9,  27,  14,   7,  27,  29,   2,   3,  18,   9,  27,  18,  12,  21,  23,  24,  11,  10,  21,  14,   7,  14,  15,   2,  20,  14,  21,  24,  22,  19,  24,  16,   9,  17,   9,  13,  17,   9,  16,  14,  29,  11,  14,   3,   8,  27,   9,  14,  24,  13,  12,   6,  32,  14,  20,  16,  21,  26,  15,  24,  22,  13,  23,  20,  16,  30,  24,  15,  24,  19,  11,  21,  26,   3,  28,  27,  20,  20,  19,  32,   8,  24,   3,   3,   0,  29,   4,   7,  16,  13,  16,   5,   1,   2,  25,   8,   7,  19,   1,  17,   7,  25,   6,  19,  14,  16,  10,   5,  22,   8,  13,  15,   6,  24,  15,  18,   4,  17,  14,   2,  18,  20,   9,  11,  20,   0,   5,  13,  24,  10,  12,   7,  12,  29,  21,  27,  23,  25,  19,   0,  26,  22,   3,  14,   6,  30,  19,  23,  17,  20,  30,  11,  26,  31,  15,  15,  19,  24,  25,   6,  20,  13,   3,  16,   3,  13,  28,  16,   4,  11,   3,  11,  15,   4,  14,  27,  22,  23,  30,  26,   1,  16,  17,  13,  12,  31,   2,  23,  12,  12,   6,   2,   5,   2,  23,   6,  18,  31,  16,  21,  15,   8,  20,  30,   7,  15,  11,  11,  26,  17,  19,  19,  12,  26,  23,   3,  25,  19,   1,   7,  16,  24,  13,   7,  16,  20,  18,  28,   8,  15,   7,  28,  13,  23,  29,  18,   4,  11,   4,  21,  16,  28,  13,  16,  15,   7,  13,  14,  20,   4,   8,  10,  19,  12,   5,  14,   4,  22,  27,  16,  23,   9,  26,  16,  19,   6,   8,  16,  32,  16,  16,  14,  31,   4,   5,  16,  11,  16,  31,   9,  21,   7,   9,  11,   8,  25,  19,   8,  22,  21,   9,  16,   2,  23,  22,  28,   6,  26,  17,  16,  15,  20,   9,  17,  26,   0,  29,  22,  22,   9,  27,   9,   7,   7,  11,  10,  15,   9,  15,  21,   5,  16,   7,   2,  13,   8,  27,  24,  22,  14,  26,  12,  10,  20,  30,   2,   9,  27,  12,  23,  28,   4,  20,   1,   9,  13,   1,  16,  27,  31,  26,  16,   7,   4,  24,   2,  27,  25,   6,  32,  10,  16,  27,  23,   1,  15,  12,   2,  27,  13,  12,   3,  29,  19,   9,  21,   7,  21,  14,   9,  12,   9,  24,  20,  19,  29,  27,  21,  18,   9,  16,  26,  17,  10,  21,  29,   8,  29,   5,  15,  15,  17,  23,  16,  18,  26,  11,  20,   4,  31,   3,  16,  26,  21,  16,  26,  21,  30,   5,  31,  15,  19,  24,  17,   1,  31,  13,  23,  24,   0,  25,  18,  18,  22,  16,  14,   2,  20,  14,   5,  16,   8,  14,  16,  24,  22,   1,   5,  11,  10,  16,   3,  17,  26,  14,  13,  18,  21,   0,  26,   4,   5,  16,  25,  21,  23,  28,  26,  14,  10,   5,  13,  20,  12,  12,  27,  20,  15,  29,  23,  19,  28,  19,  31,  29,  11,   7,   3,  16,   9,  23,  13,   4,  21,  31,  27,   2,   0,  22,   5,  22,  25,  23,  28,   5,   7,  16,  20,  10,  32,  24,  32,  26,  16,   5,  22,  24,   7,   3,  12,  31,  17,  12,  25,  19,  15,  18,  32,  19,  11,  28,  18,  24,  12,  24,  16,  13,  32,  16,   9,  10,  21,  20,  11,  32,  16,  25,   8,  32,  19,  19,   9,  15,   2,   9,   3,  31,  20,  17,  13,  13,  25,  26,  14,   1,  14,  18,   0,  19,  27,  32,   8,  23,  16,  16,  29,  22,  22,   6,  28,  26,  14,  26,  15,   8,  16,  31,  23,  25,  27,   8,  10,   0,  29,   8,  32,  19,   2,  25,  19,  21,   0,  29,  13,  27,  14,  17,   8,   0,   8,   9,  14,   1,  20,  16,  22,   4,  20,  14,   7,  28,  18,   3,  13,   8,   7,  21,  14,  13,  31,  11,  11,  22,  12,  17,  17,   6,   9,  26,  19,  20,  28,  26,  15,   7,  10,  22,  13,  19,   6,  12,  14,  12,  29,   3,  25,  22,  10,  21,  12,  24,  23,  31,  22,  27,  14,  30,  11,   9,  17,  12,  17,  11,   9,   5,  19,   0,   8,  19,  20,  31,  10,   9,  27,  23,  24,   0,  10,  21,   7,  23,  17,  11,  15,  17,  16,   8,  32,  20,  26,   6,  26,  31,   0,  19,  27,  28,  17,   7,   7,  15,  30,   9,  14,  17,  32,  31,  22,  16,  19,   7,  28,  16,  28,   4,   4,  18,  23,   4,  31,  24,  20,  10,  16,   0,  16,   9,  13,   4,  13,  10,  27,  11,  16,   0,  27,   9,  16,  29,  21,   7,  15,   3,  32,   0,  15,  29,  15,  22,  24,  16,  16,  11,  18,  17,   5,  29,  14,  16,   9,  18,  27,  15,  12,  13,  16,  29,  32,  23,  16,   0,  20,  18,  27,   6,  26,  21,   2,  21,  14,  28,  25,  17,  27,  13,  13,  18,   5,  27,  13,  24,  18,   8,  27,  16,  15,   3,   6,  22,   0,   3,   8,   7,  13,  24,  16,   6,  16,  14,  27,  13,  10,  28,  31,  19,  24,  10,  27,  25,  23,  30,  19,  16,   1,  15,  10,   1,  15,  19,  16,  28,   7,   6,  14,  11,   6,  24,  16,   4,   6,   3,  27,   4,  16,  31,   9,   9,  16,  26,  13,  17,  18,  17,  29,  20,   6,  20,  14,  27,  17,  22,  31,  23,  11,  20,  12,  31,  14,  23,  26,   4,   0,  24,  13,  13,  16,  15,  31,  14,  16,  20,   7,  27,  16,  23,  16,   6,  10,  21,   0,  30,  16,  21,  30,  24,  20,  20,   2,  15,   1,   7,   2,  23,  23,  20,   7,  16,  15,   6);
	constant test : int_vector_8bit(1023 downto 0) := (6, 15, 16, 7, 20, 23, 23, 2, 7, 1, 15, 2, 20, 20, 24, 30, 21, 16, 30, 0, 21, 10, 6, 16, 23, 16, 27, 7, 20, 16, 14, 31, 15, 16, 13, 13, 24, 0, 4, 26, 23, 14, 31, 12, 20, 11, 23, 31, 22, 17, 27, 14, 20, 6, 20, 29, 17, 18, 17, 13, 26, 16, 9, 9, 31, 16, 4, 27, 3, 6, 4, 16, 24, 6, 11, 14, 6, 7, 28, 16, 19, 15, 1, 10, 15, 1, 16, 19, 30, 23, 25, 27, 10, 24, 19, 31, 28, 10, 13, 27, 14, 16, 6, 16, 24, 13, 7, 8, 3, 0, 22, 6, 3, 15, 16, 27, 8, 18, 24, 13, 27, 5, 18, 13, 13, 27, 17, 25, 28, 14, 21, 2, 21, 26, 6, 27, 18, 20, 0, 16, 23, 32, 29, 16, 13, 12, 15, 27, 18, 9, 16, 14, 29, 5, 17, 18, 11, 16, 16, 24, 22, 15, 29, 15, 0, 32, 3, 15, 7, 21, 29, 16, 9, 27, 0, 16, 11, 27, 10, 13, 4, 13, 9, 16, 0, 16, 10, 20, 24, 31, 4, 23, 18, 4, 4, 28, 16, 28, 7, 19, 16, 22, 31, 32, 17, 14, 9, 30, 15, 7, 7, 17, 28, 27, 19, 0, 31, 26, 6, 26, 20, 32, 8, 16, 17, 15, 11, 17, 23, 7, 21, 10, 0, 24, 23, 27, 9, 10, 31, 20, 19, 8, 0, 19, 5, 9, 11, 17, 12, 17, 9, 11, 30, 14, 27, 22, 31, 23, 24, 12, 21, 10, 22, 25, 3, 29, 12, 14, 12, 6, 19, 13, 22, 10, 7, 15, 26, 28, 20, 19, 26, 9, 6, 17, 17, 12, 22, 11, 11, 31, 13, 14, 21, 7, 8, 13, 3, 18, 28, 7, 14, 20, 4, 22, 16, 20, 1, 14, 9, 8, 0, 8, 17, 14, 27, 13, 29, 0, 21, 19, 25, 2, 19, 32, 8, 29, 0, 10, 8, 27, 25, 23, 31, 16, 8, 15, 26, 14, 26, 28, 6, 22, 22, 29, 16, 16, 23, 8, 32, 27, 19, 0, 18, 14, 1, 14, 26, 25, 13, 13, 17, 20, 31, 3, 9, 2, 15, 9, 19, 19, 32, 8, 25, 16, 32, 11, 20, 21, 10, 9, 16, 32, 13, 16, 24, 12, 24, 18, 28, 11, 19, 32, 18, 15, 19, 25, 12, 17, 31, 12, 3, 7, 24, 22, 5, 16, 26, 32, 24, 32, 10, 20, 16, 7, 5, 28, 23, 25, 22, 5, 22, 0, 2, 27, 31, 21, 4, 13, 23, 9, 16, 3, 7, 11, 29, 31, 19, 28, 19, 23, 29, 15, 20, 27, 12, 12, 20, 13, 5, 10, 14, 26, 28, 23, 21, 25, 16, 5, 4, 26, 0, 21, 18, 13, 14, 26, 17, 3, 16, 10, 11, 5, 1, 22, 24, 16, 14, 8, 16, 5, 14, 20, 2, 14, 16, 22, 18, 18, 25, 0, 24, 23, 13, 31, 1, 17, 24, 19, 15, 31, 5, 30, 21, 26, 16, 21, 26, 16, 3, 31, 4, 20, 11, 26, 18, 16, 23, 17, 15, 15, 5, 29, 8, 29, 21, 10, 17, 26, 16, 9, 18, 21, 27, 29, 19, 20, 24, 9, 12, 9, 14, 21, 7, 21, 9, 19, 29, 3, 12, 13, 27, 2, 12, 15, 1, 23, 27, 16, 10, 32, 6, 25, 27, 2, 24, 4, 7, 16, 26, 31, 27, 16, 1, 13, 9, 1, 20, 4, 28, 23, 12, 27, 9, 2, 30, 20, 10, 12, 26, 14, 22, 24, 27, 8, 13, 2, 7, 16, 5, 21, 15, 9, 15, 10, 11, 7, 7, 9, 27, 9, 22, 22, 29, 0, 26, 17, 9, 20, 15, 16, 17, 26, 6, 28, 22, 23, 2, 16, 9, 21, 22, 8, 19, 25, 8, 11, 9, 7, 21, 9, 31, 16, 11, 16, 5, 4, 31, 14, 16, 16, 32, 16, 8, 6, 19, 16, 26, 9, 23, 16, 27, 22, 4, 14, 5, 12, 19, 10, 8, 4, 20, 14, 13, 7, 15, 16, 13, 28, 16, 21, 4, 11, 4, 18, 29, 23, 13, 28, 7, 15, 8, 28, 18, 20, 16, 7, 13, 24, 16, 7, 1, 19, 25, 3, 23, 26, 12, 19, 19, 17, 26, 11, 11, 15, 7, 30, 20, 8, 15, 21, 16, 31, 18, 6, 23, 2, 5, 2, 6, 12, 12, 23, 2, 31, 12, 13, 17, 16, 1, 26, 30, 23, 22, 27, 14, 4, 15, 11, 3, 11, 4, 16, 28, 13, 3, 16, 3, 13, 20, 6, 25, 24, 19, 15, 15, 31, 26, 11, 30, 20, 17, 23, 19, 30, 6, 14, 3, 22, 26, 0, 19, 25, 23, 27, 21, 29, 12, 7, 12, 10, 24, 13, 5, 0, 20, 11, 9, 20, 18, 2, 14, 17, 4, 18, 15, 24, 6, 15, 13, 8, 22, 5, 10, 16, 14, 19, 6, 25, 7, 17, 1, 19, 7, 8, 25, 2, 1, 5, 16, 13, 16, 7, 4, 29, 0, 3, 3, 24, 8, 32, 19, 20, 20, 27, 28, 3, 26, 21, 11, 19, 24, 15, 24, 30, 16, 20, 23, 13, 22, 24, 15, 26, 21, 16, 20, 14, 32, 6, 12, 13, 24, 14, 9, 27, 8, 3, 14, 11, 29, 14, 16, 9, 17, 13, 9, 17, 9, 16, 24, 19, 22, 24, 21, 14, 20, 2, 15, 14, 7, 14, 21, 10, 11, 24, 23, 21, 12, 18, 27, 9, 18, 3, 2, 29, 27, 7, 14, 27, 9, 29, 7, 15, 7, 10, 7, 7, 15, 11, 16, 22, 22, 27, 7, 6, 20, 30, 25, 16, 27, 15, 20, 13, 19, 17, 17, 17, 21, 29, 22, 6, 5, 12, 19, 7, 25, 11, 20, 16, 19, 11, 28, 20, 21, 21, 19, 18, 22, 14, 13, 26, 1, 31, 9, 15, 20, 11, 15, 20, 32, 4, 27, 27, 19, 18, 18, 24, 15, 11, 19, 14, 20, 23, 1, 20, 10, 29, 5, 15, 22, 14, 20, 5, 13, 14, 8, 27, 18, 11, 17, 10, 8, 24, 6, 9, 7, 10, 24, 17, 9, 10, 15, 16, 3, 7);
end package Amogh_pkg;
